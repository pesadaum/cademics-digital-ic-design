module sample ();

typedef enum bit [3:0] {t = 2'b2, s = 4'b4, w=3'b5} states;


endmodule